library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use STD.textio.all; -- Required for freading a file

entity instruction_memory is
	port (
		read_address: in STD_LOGIC_VECTOR (31 downto 0);
		instruction: out STD_LOGIC_VECTOR (31 downto 0)
	);
end instruction_memory;


architecture behavioral of instruction_memory is	  

    -- 128 byte instruction memory (32 rows * 4 bytes/row)
    type mem_array is array(0 to 31) of STD_LOGIC_VECTOR (31 downto 0);
    signal data_mem: mem_array := (
		  "00100000000010000000000001000010", -- addi $t0, $0, 42
		  "00001000000000000000000000001000", -- j later
		  "00100000000010010000000000000100", -- earlier: addi $t1, $0 ,4
		  "00000001000010010101000000100010", --          sub  $t2, $t0, $t1 
		  "00000001010010000101100000100101", -- 			  or $t3, $t2,$t0
		  "10101100000010110000000000101100", --          sw $t3, 2C($0)   
		  "10001101001011000000000000101000", --          lw $t4, 28($t1)
		  "00001000000000000000000000000111", -- j done              
		  "00010000000000001111111111111001", -- beq $0, $0 , earlier 
        "00000000000000000000000000000000",  
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",  
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
		  "00000000000000000000000000000000"
    );

    begin

    -- Since the registers are in multiples of 4 bytes, we can ignore the last two bits
    instruction <= data_mem(to_integer(unsigned(read_address(31 downto 2))));

end behavioral;
